module main

// TODO : Add more
fn main() {
	
}
