module main

import vmonkey

fn main() {
	lexer := vmonkey.new_lexer('test')
}
